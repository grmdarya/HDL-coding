library verilog;
use verilog.vl_types.all;
entity COMPARATOR_vlg_tst is
end COMPARATOR_vlg_tst;
